	// Calculator operation defines
  `define ADD 2'b00
  `define SUB 2'b01
  `define MUL 2'b10
  `define DIV 2'b11
  `define LOW  0
  `define HIGH 1
  `define MAX_TIME_TAKEN_BY_ONE_TRANS 1us
	`define DEFAULT_DELAY_BTWN_TXNS 		10
	`define DEFAULT_STALL_PROBABILITY 	50
//------------------------------------------------  
