package calci_pkg;
	typedef virtual calci_if calci_vif ;
	`include "calci_defines.sv"
	`include "calci_trans.sv"
	`include "calci_config.sv"
	`include "calci_gen.sv"
	`include "calci_driver.sv"
	`include "calci_sig_cov.sv"
	`include "calci_monitor.sv"
	`include "calci_ref_model.sv"
	`include "calci_trans_cov.sv"
	`include "calci_sb.sv"
	`include "calci_env.sv"
	`include "calci_test.sv"
//------------------------------------------------  
endpackage
